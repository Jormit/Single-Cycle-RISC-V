module control (
);


endmodule
